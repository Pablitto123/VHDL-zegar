----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:58:07 05/16/2021 
-- Design Name: 
-- Module Name:    zegar - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity zegar is
    Port ( 
			  Clk : in STD_LOGIC;
			  CA1 : out  STD_LOGIC;
           CB1 : out  STD_LOGIC;
           CC1 : out  STD_LOGIC;
           CD1 : out  STD_LOGIC;
			  CE1 : out  STD_LOGIC;
           CF1 : out  STD_LOGIC;
           CG1 : out  STD_LOGIC;
			  CA2 : out  STD_LOGIC;
           CB2 : out  STD_LOGIC;
           CC2 : out  STD_LOGIC;
           CD2 : out  STD_LOGIC;
			  CE2 : out  STD_LOGIC;
           CF2 : out  STD_LOGIC;
           CG2 : out  STD_LOGIC;
			  CA3 : out  STD_LOGIC;
           CB3 : out  STD_LOGIC;
           CC3 : out  STD_LOGIC;
           CD3 : out  STD_LOGIC;
			  CE3 : out  STD_LOGIC;
           CF3 : out  STD_LOGIC;
           CG3 : out  STD_LOGIC
			  );
end zegar;

architecture Behavioral of zegar is

begin


end Behavioral;

